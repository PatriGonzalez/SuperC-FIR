
* **********************************************************************
* Author      : LPGG
* Date        : 09/10/2020
* Description : Inhibit element
* Notes       :
*  - Taken from Superconducting-Temporal-Logic 
*    https://github.com/UCSBarchlab/Superconducting-Temporal-Logic.git
*  - The INHIBIT operator receives two input signals: one inhibiting and one data signal. 
*    An output pulse is emitted only if the signal arrives before the inhibiting one. 
*    To implement INHIBIT in RSFQ we use a single INVERTER. According to the INVERTER’s 
*    specification, if a data pulse arrives, the next clock pulse reads out “0”; 
*    otherwise, it reads out “1”. Thus, if we route the data signal 
*    to the inverter’s clock port and the inhibiting signal 
*    to its data port, this component will act exactly as an INHIBIT operator 
*    for our logic.
*  - The jjr element is defined at a higher level
* **********************************************************************


.subckt inhibit INH D OUT VBIAS
   X0 INH D OUT VBIAS inv
.ends inhibit


