
* **********************************************************************
* Author      : LPGG
* Date        : 09/10/2020
* Description : Simple JTL circuit element
* Notes       :
*  - Taken from Superconducting-Temporal-Logic 
*    https://github.com/UCSBarchlab/Superconducting-Temporal-Logic.git
*  - The jjr element is defined at a higher level
* **********************************************************************

.subckt jtl IN OUT VBIAS

B0 5 7 9 jjr ics=250uA
RS0 5 7 2.7
B1 6 8 10 jjr ics=250uA
RS1 6 8 2.7

LP0 7 0 .1pH
LP1 8 0 .1pH

LT0 IN 5 2.1pH
LT1 5 4 2.1pH
LT2 4 6 2.1pH
LT3 6 OUT 2.1pH

R0 VBIAS 4 29

.ends jtl

 
