
.subckt balancer IN1 IN2 OUT1 OUT2 VBIAS

X0 IN1_1 IN2_1 CLK VBIAS merge
X1 CLK s1a s1b VBIAS tff2

X2 IN1_2 s1a_0 s1b_0 c1a c2a VBIAS dff2
X3 IN2_2 s1a_1 s1b_1 c2b c1b VBIAS dff2

X4 c1a c1b clk1 VBIAS merge
X5 c2a c2b clk2 VBIAS merge
X6 IN1_3 clk1_0 clk2_0 y1a y2a VBIAS dff2
X7 IN2_3 clk2_1 clk1_1 y1b y2b VBIAS dff2

X8 y1a y1b OUT1 VBIAS merge
X9 y2a y2b OUT2 VBIAS merge

*- Spliting
X10 IN1   IN1_0 IN1_1  VBIAS split
X11 IN1_0 IN1_2 IN1_3  VBIAS split
X12 IN2   IN2_0 IN2_1  VBIAS split
X13 IN2_0 IN2_2 IN2_3  VBIAS split
X14 s1a s1a_0 s1a_1    VBIAS split
X15 s1b s1b_0 s1b_1    VBIAS split
X16 clk1 clk1_0 clk1_1 VBIAS split
X17 clk2 clk2_0 clk2_1 VBIAS split


.ends balancer

*plot v(nT0) v(nT1) v(Set1c.Xf87) v(Set2d.Xf87) v(Set2c.Xf87) v(Set1d.Xf87) v(IN1_5j_0_del.Xf87) v(IN2_5j_0_del.Xf87) v(Q1a.Xf87) v(Q2a.Xf87) v(Q1b.Xf87) v(Q2b.Xf87)  

*plot v(nT0) v(nT1) v(Set1c.Xf87) v(Set1d.Xf87) v(Set2c.Xf87) v(nY00) v(nY01) 
*plot v(nT0) v(nT1) v(nY00) v(nY01) v(Set1c.Xf87) v(Set1d.Xf87) v(Set2c.Xf87) v(Set2d.Xf87) 
*plot v(nT0) v(nT1) v(Set1c.Xf87) v(Rst1a.Xf87) v(IN1_5j_0_del.Xf87) v(Q1a.Xf87) 
*plot v(nT0) v(nT1) v(Set2d.Xf87) v(Rst2a.Xf87) v(IN1_5j_1_del.Xf87) v(Q2a.Xf87) 
*plot v(nT0) v(nT1) v(Set2c.Xf87) v(Rst2b.Xf87) v(IN2_5j_0_del.Xf87) v(Q1b.Xf87) 
*plot v(nT0) v(nT1) v(Set1d.Xf87) v(Rst1b.Xf87) v(IN2_5j_1_del.Xf87) v(Q2b.Xf87)

*X0  IN1   IN1_0 IN1_1 VBIAS split
*X0a IN1_0 IN1_2 IN1_3 VBIAS split
*X0b IN1_2 IN1_4 IN1_5 VBIAS split
*
*X1  IN2   IN2_0 IN2_1 VBIAS split
*X1a IN2_0 IN2_2 IN2_3 VBIAS split
*X1b IN2_2 IN2_4 IN2_5 VBIAS split
*
*X3 IN2_3 IN1_3 S1 VBIAS inv
*X2 IN1_1 IN2_1 S2 VBIAS inv 
*
*X4 S1 S1a S1b VBIAS tff2
*X5 S2 S2a S2b VBIAS tff2
*
*X6 S1a S2b S3 VBIAS merge
*X7 S1b S2a S4 VBIAS merge
*
*X100 S3 Rst2 Set1_0 VBIAS split
*X101 S4 Rst1 Set2_0 VBIAS split
*
*X102 Set1_0 Set1_1 VBIAS jtl
*X103 Set1_1 Set1   VBIAS jtl
*X104 Set2_0 Set2_1 VBIAS jtl
*X105 Set2_1 Set2   VBIAS jtl
*
*X108 Set1  Set1a Set1b VBIAS split 
*X108a Set1a Set1c Set1d VBIAS split
*
*X109 Set2  Set2a Set2b VBIAS split 
*X109a Set2a Set2c Set2d VBIAS split 
*
*X110 Rst1 Rst1a Rst1b VBIAS split 
*X111 Rst2 Rst2a Rst2b VBIAS split 
*
*X8a IN1_5  IN1_5a VBIAS jtl
*X8b IN1_5a IN1_5b VBIAS jtl
*X8c IN1_5b IN1_5c VBIAS jtl
*X8d IN1_5c IN1_5d VBIAS jtl
*X8e IN1_5d IN1_5e VBIAS jtl
*X8f IN1_5e IN1_5f VBIAS jtl
*X8g IN1_5f IN1_5g VBIAS jtl
*X8h IN1_5g IN1_5h VBIAS jtl
*X8i IN1_5h IN1_5i VBIAS jtl
*X8j IN1_5i IN1_5j VBIAS jtl
*X8o IN1_5j IN1_5j_0 IN1_5j_1 VBIAS split
*X8ja IN1_5j_0 IN1_5j_0_del VBIAS jtl
*X8jb IN1_5j_1 IN1_5j_1_del VBIAS jtl
*
*
*X9a IN2_5  IN2_5a VBIAS jtl
*X9b IN2_5a IN2_5b VBIAS jtl
*X9c IN2_5b IN2_5c VBIAS jtl
*X9d IN2_5c IN2_5d VBIAS jtl
*X9e IN2_5d IN2_5e VBIAS jtl
*X9f IN2_5e IN2_5f VBIAS jtl
*X9g IN2_5f IN2_5g VBIAS jtl
*X9h IN2_5g IN2_5h VBIAS jtl
*X9i IN2_5h IN2_5i VBIAS jtl
*X9j IN2_5i IN2_5j VBIAS jtl
*X9o IN2_5j IN2_5j_0 IN2_5j_1 VBIAS split
*X9ja IN2_5j_0 IN2_5j_0_del VBIAS jtl
*X9jb IN2_5j_1 IN2_5j_1_del VBIAS jtl
*
*X8 Set1c NC0 Rst1a IN1_5j_0_del Q1a VBIAS ndro_il
*X9 Set2d NC1 Rst2a IN1_5j_1_del Q2a VBIAS ndro_il
*
*
*X10 Set2c NC2 Rst2b IN2_5j_0_del Q1b VBIAS ndro_il
*X11 Set1d NC3 Rst1b IN2_5j_1_del Q2b VBIAS ndro_il
*
*X16 Q1a Q1b OUT1 VBIAS merge
*X18 Q2a Q2b OUT2 VBIAS merge
