
* **********************************************************************
* Author      : LPGG
* Date        : 09/10/2020
* Description : 2 outputs Toggle flipflop
* Notes       :
*  - Implemented by Meriam Bautista (mgbautista@lbl.gov)
*  - The jjr element is defined at a higher level
* **********************************************************************


.subckt tff2 IN OUT1 OUT2 VBIAS

B1  1 0 n1 jjr ics=125uA
RS1 1 0 5.4

B2  2 0 n2 jjr ics=192uA
RS2 2 0 3.5

*B3  1 3 n3 jjr ics=302uA
*RS3 1 3 0.4

*B3  1 3 n3 jjr ics=250uA
*RS3 1 3 2.7

B3  1 3 n3 jjr ics=200uA
RS3 1 3 3.2

B4  2 4 n4 jjr ics=125uA
RS4 2 4 5.4

B5  5 0 n5 jjr ics=250uA
RS5 5 0 2.7

B6  6 0 n6 jjr ics=250uA
RS6 6 0 2.7

B7  7 0 n7 jjr ics=125uA
RS7 7 0 5.4

B8  8 0 n8 jjr ics=192uA
RS8 8 0 3.5

B9  9 0 n9 jjr ics=192uA
RS9 9 0 3.5

B10  10 0 n10 jjr ics=250uA
RS10 10 0 2.7

L1   1    2 8.00pH
L2   3   12 0.14pH
L3  12    4 1.87pH
L4  IN    5 2.67pH
L5   5   11 1.33pH
L6  11    6 0.80pH
L7   6   12 0.27pH
L8   1    7 8.00pH
L9   7   14 4.00pH
L10 14    8 1.33pH
L11  8 OUT1 4.00pH
L12  2    9 5.33pH
L13  9   13 4.00pH
L14 13   10 1.33pH
L15 10 OUT2 4.00pH


*R1 VBIAS 11 22
*R2 VBIAS 13 32
*R3 VBIAS 14 39

R1 VBIAS 11 20
R2 VBIAS 13 37
R3 VBIAS 14 32

.ends tff2
