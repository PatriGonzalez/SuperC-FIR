
******************************
* Specify simulation options
******************************
.tran 0.5p 17662.24p
*.tran 0.5p 500p
.options maxdata=3500000

******************************
* Specity Inputs
******************************
V0 VCC 0 pwl 0 0 10p 10m

*- INFO: Used to SET the coefficient NDROs
V1 1 0 pulse 0 50m 50p 50p 10p 10p 1m
R1 1 2 100
X1_sfq 2 SET_COEF VCC dcsfq

*- INFO: Used to RESET the coefficient NDROs
V2 3 0 pulse 0 0 0p 50p 10p 10p 1900p
R2 3 4 100
X2_sfq 4 RST_COEF VCC dcsfq

*- INFO: Used to SET the multipliers
V3 5 0 pulse 0 50m 224p 50p 10p 10p 1m
R3 5 6 100
X3_sfq 6 INIT VCC dcsfq

*- INFO: No VCO, just an external CLK with delay 10p
V4 7 0 pulse 0 50m 10p 50p 10p 10p 128.32p
R4 7 8 100
X4_sfq 8 CLK VCC dcsfq

******************************
* Circuit 
******************************
  Xf0 CLK CLKa0 CLKa VCC split
  Xf1 CLKa0 CLKb0 CLKb VCC split
  Xf2 CLKb0 CLKc0 CLKc VCC split
  Xf3 CLKc0 CLKd0 CLKd VCC split

  Xf4 INIT RST_EPOCHa INIT_M VCC merge
  Xf5 INIT_M INIT_Ma SET_EPOCH VCC split
  Xf6 INIT_Ma INIT0 CLKa VCC dff_il
  Xf7 INIT0 INIT0a INIT0b VCC split
  Xf8 INIT0a INIT1 CLKc VCC dff_il
  Xf9 INIT1 NC0 RST_EPOCHd CLKd CLK_Mult0 VCC ndro_il
  Xf10 CLK_Mult0 CLK_Mult VCC jtl
  Xf11 INIT0b NC1 RST_EPOCHc CLKb CLK_Gen0 VCC ndro_il
  Xf12 CLK_Gen0 CLK_Gen VCC jtl

  Xf13 nP6 RST_EPOCHb RST_EPOCHe VCC split
  Xf14 RST_EPOCHb RST_EPOCHc RST_EPOCHd VCC split
  Xf15 RST_EPOCHe RST_EPOCHa RST_EPOCH VCC split

*INFO: Instantiate toggle flipflops
  Xf16 CLK_Gen nP0a nP0 VCC tff2
  Xf17 nP0 nP1a nP1 VCC tff2
  Xf18 nP1 nP2a nP2 VCC tff2
  Xf19 nP2 nP3a nP3 VCC tff2
  Xf20 nP3 nP4a nP4 VCC tff2
  Xf21 nP4 nP5a nP5 VCC tff2
  Xf22 nP5 nP6a nP6 VCC tff2

*- INFO: Merge the pulses
  Xf23 n00 nArm0 VCC merge_arm 
  Xf24 n01 nArm0 VCC merge_arm 
  Xf25 n02 nArm0 VCC merge_arm 
  Xf26 n03 nArm0 VCC merge_arm 
  Xf27 n04 nArm0 VCC merge_arm 
  Xf28 n05 nArm0 VCC merge_arm 
  Xf29 n06 nArm0 VCC merge_arm 
  B30 30_11 30_13 30_19 jjr ics=250uA
  RS30 30_11 30_13 2.7
  L30_1 30_5 30_11   2.6pH
  L30_2 30_11 nCoef0 2pH
  LP30_3 nArm0 30_5 .2pH
  LP30_5 30_13 0 .03pH

  Xf30 n10 nArm1 VCC merge_arm 
  Xf31 n11 nArm1 VCC merge_arm 
  Xf32 n12 nArm1 VCC merge_arm 
  Xf33 n13 nArm1 VCC merge_arm 
  Xf34 n14 nArm1 VCC merge_arm 
  Xf35 n15 nArm1 VCC merge_arm 
  Xf36 n16 nArm1 VCC merge_arm 
  B37 37_11 37_13 37_19 jjr ics=250uA
  RS37 37_11 37_13 2.7
  L37_1 37_5 37_11   2.6pH
  L37_2 37_11 nCoef1 2pH
  LP37_3 nArm1 37_5 .2pH
  LP37_5 37_13 0 .03pH

  Xf37 n20 nArm2 VCC merge_arm 
  Xf38 n21 nArm2 VCC merge_arm 
  Xf39 n22 nArm2 VCC merge_arm 
  Xf40 n23 nArm2 VCC merge_arm 
  Xf41 n24 nArm2 VCC merge_arm 
  Xf42 n25 nArm2 VCC merge_arm 
  Xf43 n26 nArm2 VCC merge_arm 
  B44 44_11 44_13 44_19 jjr ics=250uA
  RS44 44_11 44_13 2.7
  L44_1 44_5 44_11   2.6pH
  L44_2 44_11 nCoef2 2pH
  LP44_3 nArm2 44_5 .2pH
  LP44_5 44_13 0 .03pH

  Xf44 n30 nArm3 VCC merge_arm 
  Xf45 n31 nArm3 VCC merge_arm 
  Xf46 n32 nArm3 VCC merge_arm 
  Xf47 n33 nArm3 VCC merge_arm 
  Xf48 n34 nArm3 VCC merge_arm 
  Xf49 n35 nArm3 VCC merge_arm 
  Xf50 n36 nArm3 VCC merge_arm 
  B51 51_11 51_13 51_19 jjr ics=250uA
  RS51 51_11 51_13 2.7
  L51_1 51_5 51_11   2.6pH
  L51_2 51_11 nCoef3 2pH
  LP51_3 nArm3 51_5 .2pH
  LP51_5 51_13 0 .03pH


*- INFO: Now the multipliers
  Xf51 CLK_Mult CLK0s CLK0 VCC split
  Xf52 nCoef0 nCoef0a nCoef0b VCC split
  Xf53 nCoef0b CLK0 nCoef0c VCC inv
  Xf54 nX0 nX0a nX0b VCC split
  Xf55 SET_EPOCH SET_EPOCH0s SET_EPOCH0 VCC split
  Xf56 RST_EPOCH RST_EPOCH0s RST_EPOCH0 VCC split
  Xf57 SET_EPOCH0 NC0a nX0a nCoef0a nT0a VCC ndro_il
  Xf58 nX0b NC0b RST_EPOCH0 nCoef0c nT0b VCC ndro_il
  Xf59 nT0a nT0b nT0 VCC merge

  Xf60 CLK0s CLK1s CLK1 VCC split
  Xf61 nCoef1 nCoef1a nCoef1b VCC split
  Xf62 nCoef1b CLK1 nCoef1c VCC inv
  Xf63 nX1 nX1a nX1b VCC split
  Xf64 SET_EPOCH0s SET_EPOCH1s SET_EPOCH1 VCC split
  Xf65 RST_EPOCH0s RST_EPOCH1s RST_EPOCH1 VCC split
  Xf66 SET_EPOCH1 NC1a nX1a nCoef1a nT1a VCC ndro_il
  Xf67 nX1b NC1b RST_EPOCH1 nCoef1c nT1b VCC ndro_il
  Xf68 nT1a nT1b nT1 VCC merge

  Xf69 CLK1s CLK2s CLK2 VCC split
  Xf70 nCoef2 nCoef2a nCoef2b VCC split
  Xf71 nCoef2b CLK2 nCoef2c VCC inv
  Xf72 nX2 nX2a nX2b VCC split
  Xf73 SET_EPOCH1s SET_EPOCH2s SET_EPOCH2 VCC split
  Xf74 RST_EPOCH1s RST_EPOCH2s RST_EPOCH2 VCC split
  Xf75 SET_EPOCH2 NC2a nX2a nCoef2a nT2a VCC ndro_il
  Xf76 nX2b NC2b RST_EPOCH2 nCoef2c nT2b VCC ndro_il
  Xf77 nT2a nT2b nT2 VCC merge

  Xf78 CLK2s CLK3s CLK3 VCC split
  Xf79 nCoef3 nCoef3a nCoef3b VCC split
  Xf80 nCoef3b CLK3 nCoef3c VCC inv
  Xf81 nX3 nX3a nX3b VCC split
  Xf82 SET_EPOCH2s SET_EPOCH3s SET_EPOCH3 VCC split
  Xf83 RST_EPOCH2s RST_EPOCH3s RST_EPOCH3 VCC split
  Xf84 SET_EPOCH3 NC3a nX3a nCoef3a nT3a VCC ndro_il
  Xf85 nX3b NC3b RST_EPOCH3 nCoef3c nT3b VCC ndro_il
  Xf86 nT3a nT3b nT3 VCC merge


*- INFO: Now the Adder
  Xf87 nT0 nT1 nY00 nY01 VCC balancer
  Xf88 nT2 nT3 nY02 nY03 VCC balancer

  Xf89 nY00 nY02d nY10 nY11a VCC balancer

  Xf90 nY11a nY11 VCC jtl  

  X1004 nY02 nY02d VCC jtl
  *X1005 nY02d_0 nY02d VCC jtl
  *X1006 nY02d_1 nY02d VCC jtl

